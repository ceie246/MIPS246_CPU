library verilog;
use verilog.vl_types.all;
entity top_vga_tb is
end top_vga_tb;
