library verilog;
use verilog.vl_types.all;
entity top_core_tb is
end top_core_tb;
