library verilog;
use verilog.vl_types.all;
entity top_itype_tb is
end top_itype_tb;
