library verilog;
use verilog.vl_types.all;
entity wram2asciiram_addr_tb is
end wram2asciiram_addr_tb;
