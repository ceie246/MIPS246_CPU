library verilog;
use verilog.vl_types.all;
entity kb2ascii is
    generic(
        ascii_1         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1);
        ascii_2         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        ascii_3         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1);
        ascii_4         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        ascii_5         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1);
        ascii_6         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0);
        ascii_7         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1);
        ascii_8         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0);
        ascii_9         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1);
        ascii_0         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        ascii_a         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        ascii_b         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0);
        ascii_c         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        ascii_d         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        ascii_e         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1);
        ascii_f         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        ascii_g         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        ascii_h         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        ascii_i         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1);
        ascii_j         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0);
        ascii_k         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1);
        ascii_l         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0);
        ascii_m         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1);
        ascii_n         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0);
        ascii_o         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1);
        ascii_p         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        ascii_q         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1);
        ascii_r         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        ascii_s         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1);
        ascii_t         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        ascii_u         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1);
        ascii_v         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0);
        ascii_w         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1);
        ascii_x         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0);
        ascii_y         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1);
        ascii_z         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0);
        ascii_wave      : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        ascii_sub       : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1);
        ascii_add       : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1);
        ascii_left_bracket: vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1);
        ascii_right_bracket: vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1);
        ascii_or        : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        ascii_colon     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1);
        ascii_quotes    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        ascii_comma     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0);
        ascii_dot       : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0);
        ascii_div       : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1);
        ascii_shift_1   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        ascii_shift_2   : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ascii_shift_3   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        ascii_shift_4   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        ascii_shift_5   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1);
        ascii_shift_6   : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        ascii_shift_7   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        ascii_shift_8   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0);
        ascii_shift_9   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        ascii_shift_0   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1);
        ascii_shift_wave: vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0);
        ascii_shift_sub : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1);
        ascii_shift_add : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1);
        ascii_shift_left_bracket: vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1);
        ascii_shift_right_bracket: vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1);
        ascii_shift_or  : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        ascii_shift_colon: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0);
        ascii_shift_quotes: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0);
        ascii_shift_comma: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        ascii_shift_dot : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0);
        ascii_shift_div : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        kb_1            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0);
        kb_2            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        kb_3            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        kb_4            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1);
        kb_5            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0);
        kb_6            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0);
        kb_7            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1);
        kb_8            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0);
        kb_9            : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        kb_0            : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        kb_a            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        kb_b            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        kb_c            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        kb_d            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        kb_e            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        kb_f            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1);
        kb_g            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        kb_h            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1);
        kb_i            : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        kb_j            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1);
        kb_k            : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        kb_l            : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1);
        kb_m            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0);
        kb_n            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1);
        kb_o            : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        kb_p            : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        kb_q            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        kb_r            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1);
        kb_s            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1);
        kb_t            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0);
        kb_u            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        kb_v            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0);
        kb_w            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1);
        kb_x            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0);
        kb_y            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1);
        kb_z            : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0);
        kb_wave         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0);
        kb_sub          : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0);
        kb_add          : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        kb_left_bracket : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        kb_right_bracket: vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1);
        kb_or           : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1);
        kb_colon        : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        kb_quotes       : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0);
        kb_comma        : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        kb_dot          : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        kb_div          : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        kb_ESC          : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0);
        kb_F1           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        kb_F2           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        kb_F3           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        kb_F4           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        kb_F5           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        kb_F6           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1);
        kb_F7           : vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        kb_F8           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        kb_F9           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        kb_F10          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        kb_F11          : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0);
        kb_F12          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        kb_TAB          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        kb_CAPS         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        kb_SHIFT_LEFT   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0);
        kb_SHIFT_RIGHT  : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        kb_CTRL         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        kb_ALT          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1);
        kb_SPACE        : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1);
        kb_ENTER        : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0);
        kb_BACK         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        kb_UP           : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1);
        kb_DOWN         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        kb_LEFT         : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1);
        kb_RIGHT        : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0)
    );
    port(
        data_in         : in     vl_logic_vector(7 downto 0);
        data_out        : out    vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ascii_1 : constant is 1;
    attribute mti_svvh_generic_type of ascii_2 : constant is 1;
    attribute mti_svvh_generic_type of ascii_3 : constant is 1;
    attribute mti_svvh_generic_type of ascii_4 : constant is 1;
    attribute mti_svvh_generic_type of ascii_5 : constant is 1;
    attribute mti_svvh_generic_type of ascii_6 : constant is 1;
    attribute mti_svvh_generic_type of ascii_7 : constant is 1;
    attribute mti_svvh_generic_type of ascii_8 : constant is 1;
    attribute mti_svvh_generic_type of ascii_9 : constant is 1;
    attribute mti_svvh_generic_type of ascii_0 : constant is 1;
    attribute mti_svvh_generic_type of ascii_a : constant is 1;
    attribute mti_svvh_generic_type of ascii_b : constant is 1;
    attribute mti_svvh_generic_type of ascii_c : constant is 1;
    attribute mti_svvh_generic_type of ascii_d : constant is 1;
    attribute mti_svvh_generic_type of ascii_e : constant is 1;
    attribute mti_svvh_generic_type of ascii_f : constant is 1;
    attribute mti_svvh_generic_type of ascii_g : constant is 1;
    attribute mti_svvh_generic_type of ascii_h : constant is 1;
    attribute mti_svvh_generic_type of ascii_i : constant is 1;
    attribute mti_svvh_generic_type of ascii_j : constant is 1;
    attribute mti_svvh_generic_type of ascii_k : constant is 1;
    attribute mti_svvh_generic_type of ascii_l : constant is 1;
    attribute mti_svvh_generic_type of ascii_m : constant is 1;
    attribute mti_svvh_generic_type of ascii_n : constant is 1;
    attribute mti_svvh_generic_type of ascii_o : constant is 1;
    attribute mti_svvh_generic_type of ascii_p : constant is 1;
    attribute mti_svvh_generic_type of ascii_q : constant is 1;
    attribute mti_svvh_generic_type of ascii_r : constant is 1;
    attribute mti_svvh_generic_type of ascii_s : constant is 1;
    attribute mti_svvh_generic_type of ascii_t : constant is 1;
    attribute mti_svvh_generic_type of ascii_u : constant is 1;
    attribute mti_svvh_generic_type of ascii_v : constant is 1;
    attribute mti_svvh_generic_type of ascii_w : constant is 1;
    attribute mti_svvh_generic_type of ascii_x : constant is 1;
    attribute mti_svvh_generic_type of ascii_y : constant is 1;
    attribute mti_svvh_generic_type of ascii_z : constant is 1;
    attribute mti_svvh_generic_type of ascii_wave : constant is 1;
    attribute mti_svvh_generic_type of ascii_sub : constant is 1;
    attribute mti_svvh_generic_type of ascii_add : constant is 1;
    attribute mti_svvh_generic_type of ascii_left_bracket : constant is 1;
    attribute mti_svvh_generic_type of ascii_right_bracket : constant is 1;
    attribute mti_svvh_generic_type of ascii_or : constant is 1;
    attribute mti_svvh_generic_type of ascii_colon : constant is 1;
    attribute mti_svvh_generic_type of ascii_quotes : constant is 1;
    attribute mti_svvh_generic_type of ascii_comma : constant is 1;
    attribute mti_svvh_generic_type of ascii_dot : constant is 1;
    attribute mti_svvh_generic_type of ascii_div : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_1 : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_2 : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_3 : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_4 : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_5 : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_6 : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_7 : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_8 : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_9 : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_0 : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_wave : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_sub : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_add : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_left_bracket : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_right_bracket : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_or : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_colon : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_quotes : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_comma : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_dot : constant is 1;
    attribute mti_svvh_generic_type of ascii_shift_div : constant is 1;
    attribute mti_svvh_generic_type of kb_1 : constant is 1;
    attribute mti_svvh_generic_type of kb_2 : constant is 1;
    attribute mti_svvh_generic_type of kb_3 : constant is 1;
    attribute mti_svvh_generic_type of kb_4 : constant is 1;
    attribute mti_svvh_generic_type of kb_5 : constant is 1;
    attribute mti_svvh_generic_type of kb_6 : constant is 1;
    attribute mti_svvh_generic_type of kb_7 : constant is 1;
    attribute mti_svvh_generic_type of kb_8 : constant is 1;
    attribute mti_svvh_generic_type of kb_9 : constant is 1;
    attribute mti_svvh_generic_type of kb_0 : constant is 1;
    attribute mti_svvh_generic_type of kb_a : constant is 1;
    attribute mti_svvh_generic_type of kb_b : constant is 1;
    attribute mti_svvh_generic_type of kb_c : constant is 1;
    attribute mti_svvh_generic_type of kb_d : constant is 1;
    attribute mti_svvh_generic_type of kb_e : constant is 1;
    attribute mti_svvh_generic_type of kb_f : constant is 1;
    attribute mti_svvh_generic_type of kb_g : constant is 1;
    attribute mti_svvh_generic_type of kb_h : constant is 1;
    attribute mti_svvh_generic_type of kb_i : constant is 1;
    attribute mti_svvh_generic_type of kb_j : constant is 1;
    attribute mti_svvh_generic_type of kb_k : constant is 1;
    attribute mti_svvh_generic_type of kb_l : constant is 1;
    attribute mti_svvh_generic_type of kb_m : constant is 1;
    attribute mti_svvh_generic_type of kb_n : constant is 1;
    attribute mti_svvh_generic_type of kb_o : constant is 1;
    attribute mti_svvh_generic_type of kb_p : constant is 1;
    attribute mti_svvh_generic_type of kb_q : constant is 1;
    attribute mti_svvh_generic_type of kb_r : constant is 1;
    attribute mti_svvh_generic_type of kb_s : constant is 1;
    attribute mti_svvh_generic_type of kb_t : constant is 1;
    attribute mti_svvh_generic_type of kb_u : constant is 1;
    attribute mti_svvh_generic_type of kb_v : constant is 1;
    attribute mti_svvh_generic_type of kb_w : constant is 1;
    attribute mti_svvh_generic_type of kb_x : constant is 1;
    attribute mti_svvh_generic_type of kb_y : constant is 1;
    attribute mti_svvh_generic_type of kb_z : constant is 1;
    attribute mti_svvh_generic_type of kb_wave : constant is 1;
    attribute mti_svvh_generic_type of kb_sub : constant is 1;
    attribute mti_svvh_generic_type of kb_add : constant is 1;
    attribute mti_svvh_generic_type of kb_left_bracket : constant is 1;
    attribute mti_svvh_generic_type of kb_right_bracket : constant is 1;
    attribute mti_svvh_generic_type of kb_or : constant is 1;
    attribute mti_svvh_generic_type of kb_colon : constant is 1;
    attribute mti_svvh_generic_type of kb_quotes : constant is 1;
    attribute mti_svvh_generic_type of kb_comma : constant is 1;
    attribute mti_svvh_generic_type of kb_dot : constant is 1;
    attribute mti_svvh_generic_type of kb_div : constant is 1;
    attribute mti_svvh_generic_type of kb_ESC : constant is 1;
    attribute mti_svvh_generic_type of kb_F1 : constant is 1;
    attribute mti_svvh_generic_type of kb_F2 : constant is 1;
    attribute mti_svvh_generic_type of kb_F3 : constant is 1;
    attribute mti_svvh_generic_type of kb_F4 : constant is 1;
    attribute mti_svvh_generic_type of kb_F5 : constant is 1;
    attribute mti_svvh_generic_type of kb_F6 : constant is 1;
    attribute mti_svvh_generic_type of kb_F7 : constant is 1;
    attribute mti_svvh_generic_type of kb_F8 : constant is 1;
    attribute mti_svvh_generic_type of kb_F9 : constant is 1;
    attribute mti_svvh_generic_type of kb_F10 : constant is 1;
    attribute mti_svvh_generic_type of kb_F11 : constant is 1;
    attribute mti_svvh_generic_type of kb_F12 : constant is 1;
    attribute mti_svvh_generic_type of kb_TAB : constant is 1;
    attribute mti_svvh_generic_type of kb_CAPS : constant is 1;
    attribute mti_svvh_generic_type of kb_SHIFT_LEFT : constant is 1;
    attribute mti_svvh_generic_type of kb_SHIFT_RIGHT : constant is 1;
    attribute mti_svvh_generic_type of kb_CTRL : constant is 1;
    attribute mti_svvh_generic_type of kb_ALT : constant is 1;
    attribute mti_svvh_generic_type of kb_SPACE : constant is 1;
    attribute mti_svvh_generic_type of kb_ENTER : constant is 1;
    attribute mti_svvh_generic_type of kb_BACK : constant is 1;
    attribute mti_svvh_generic_type of kb_UP : constant is 1;
    attribute mti_svvh_generic_type of kb_DOWN : constant is 1;
    attribute mti_svvh_generic_type of kb_LEFT : constant is 1;
    attribute mti_svvh_generic_type of kb_RIGHT : constant is 1;
end kb2ascii;
