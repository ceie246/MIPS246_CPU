library verilog;
use verilog.vl_types.all;
entity clkdiv_init_tb is
end clkdiv_init_tb;
