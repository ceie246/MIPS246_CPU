library verilog;
use verilog.vl_types.all;
entity CLK_MANAGER_tb is
end CLK_MANAGER_tb;
