`timescale 1ns / 1ps
`include "define.v"
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:50:06 09/09/2013 
// Design Name: 
// Module Name:    wram2asciiram_addr 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module wram2asciiram_addr(
		input [31:0] addr_in,
		output [`RAM_ADDR - 1:0] addr_out
    );

always @(*) begin

end

endmodule
