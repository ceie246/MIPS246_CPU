library verilog;
use verilog.vl_types.all;
entity file_write_regfiles is
    port(
        clk             : in     vl_logic;
        regfiles0       : in     vl_logic_vector(31 downto 0);
        regfiles1       : in     vl_logic_vector(31 downto 0);
        regfiles2       : in     vl_logic_vector(31 downto 0);
        regfiles3       : in     vl_logic_vector(31 downto 0);
        regfiles4       : in     vl_logic_vector(31 downto 0);
        regfiles5       : in     vl_logic_vector(31 downto 0);
        regfiles6       : in     vl_logic_vector(31 downto 0);
        regfiles7       : in     vl_logic_vector(31 downto 0);
        regfiles8       : in     vl_logic_vector(31 downto 0);
        regfiles9       : in     vl_logic_vector(31 downto 0);
        regfiles10      : in     vl_logic_vector(31 downto 0);
        regfiles11      : in     vl_logic_vector(31 downto 0);
        regfiles12      : in     vl_logic_vector(31 downto 0);
        regfiles13      : in     vl_logic_vector(31 downto 0);
        regfiles14      : in     vl_logic_vector(31 downto 0);
        regfiles15      : in     vl_logic_vector(31 downto 0);
        regfiles16      : in     vl_logic_vector(31 downto 0);
        regfiles17      : in     vl_logic_vector(31 downto 0);
        regfiles18      : in     vl_logic_vector(31 downto 0);
        regfiles19      : in     vl_logic_vector(31 downto 0);
        regfiles20      : in     vl_logic_vector(31 downto 0);
        regfiles21      : in     vl_logic_vector(31 downto 0);
        regfiles22      : in     vl_logic_vector(31 downto 0);
        regfiles23      : in     vl_logic_vector(31 downto 0);
        regfiles24      : in     vl_logic_vector(31 downto 0);
        regfiles25      : in     vl_logic_vector(31 downto 0);
        regfiles26      : in     vl_logic_vector(31 downto 0);
        regfiles27      : in     vl_logic_vector(31 downto 0);
        regfiles28      : in     vl_logic_vector(31 downto 0);
        regfiles29      : in     vl_logic_vector(31 downto 0);
        regfiles30      : in     vl_logic_vector(31 downto 0);
        regfiles31      : in     vl_logic_vector(31 downto 0)
    );
end file_write_regfiles;
