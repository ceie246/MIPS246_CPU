library verilog;
use verilog.vl_types.all;
entity file_write_tb is
end file_write_tb;
