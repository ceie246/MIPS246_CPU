library verilog;
use verilog.vl_types.all;
entity state_machine_tb is
end state_machine_tb;
