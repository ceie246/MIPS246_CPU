library verilog;
use verilog.vl_types.all;
entity segmentcu_tb is
end segmentcu_tb;
