`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:45:52 06/10/2013 
// Design Name: 
// Module Name:    FEPU 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module FEPU(
		input clk,
		input rst,
		output [31:0] FEPU_BEPU_select, //lw����swƬѡ�ź�
		output FEPU_BEPU_w, //дmemory��IO�ź�
		output [31:0] FEPU_BEPU_data, //֮������inout
		output [31:0] FEPU_BEPU_addr
    );

wire [31:0] bc_cpu_data, cpu_bc_data;
wire [31:0] cpu_bc_addr;
wire cpu_bc_rw;

top_cpu cpu(clk, rst, bc_cpu_data, cpu_bc_data, cpu_bc_addr, cpu_bc_w);
bus_controller bc(cpu_bc_addr, cpu_bc_w, FEPU_BEPU_select, FEPU_BEPU_w);//FEPU_BEPU_data,

assign FEPU_BEPU_addr = 32'b0;
assign bc_cpu_data = 32'b0;
assign FEPU_BEPU_data = cpu_bc_data;

endmodule
